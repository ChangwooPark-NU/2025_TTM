`timescale 1ns/1ps 

module regfile2 ( 
	input logic clk, 
	input logic [6:0] a1, a2, a3, a4,
	output logic [127:0] bias
); 
	logic [31:0] mem [0:127] = '{ 
		32'hFFFFFCA3,
		32'hFFFFFA81,
		32'h000000CF,
		32'h0000014C,
		32'hFFFFFE8B,
		32'h00000303,
		32'hFFFFFF9C,
		32'h000001B9,
		32'h00000577,
		32'h00000543,
		32'h0000047F,
		32'hFFFFFDAC,
		32'h0000001F,
		32'hFFFFFE4F,
		32'h0000019F,
		32'h0000034E,
		32'h000000EF,
		32'hFFFFFE31,
		32'h000000F2,
		32'hFFFFFBD7,
		32'hFFFFFB15,
		32'hFFFFFF07,
		32'hFFFFFF7C,
		32'hFFFFFED1,
		32'h0000028A,
		32'h000001C6,
		32'h00000159,
		32'h00000165,
		32'hFFFFFFAE,
		32'h0000010D,
		32'hFFFFFC27,
		32'hFFFFFC6B,
		32'h000000A8,
		32'h00000386,
		32'h0000003F,
		32'h0000051E,
		32'h0000048A,
		32'hFFFFFA63,
		32'hFFFFFD69,
		32'h000001F4,
		32'hFFFFFFBB,
		32'h000001E3,
		32'hFFFFFCEA,
		32'h00000300,
		32'hFFFFFCC5,
		32'h00000062,
		32'hFFFFFB83,
		32'hFFFFFE62,
		32'h00000397,
		32'h000002E9,
		32'hFFFFFBF2,
		32'h00000338,
		32'hFFFFFF2C,
		32'hFFFFFBAF,
		32'h00000519,
		32'h000001E8,
		32'h00000098,
		32'h000001C9,
		32'h0000027D,
		32'hFFFFFAEF,
		32'h00000336,
		32'h0000041B,
		32'h000000B1,
		32'hFFFFFE67,
		32'h000000CB,
		32'h00000063,
		32'h000000F3,
		32'hFFFFFC82,
		32'h0000038E,
		32'h00000058,
		32'h00000055,
		32'hFFFFFDEC,
		32'h000004DF,
		32'hFFFFFBF9,
		32'hFFFFFE19,
		32'hFFFFFC35,
		32'h00000437,
		32'hFFFFFDBF,
		32'h00000019,
		32'hFFFFFF9C,
		32'h0000043E,
		32'hFFFFFB3E,
		32'hFFFFFD1B,
		32'hFFFFFA89,
		32'hFFFFFEC8,
		32'hFFFFFB27,
		32'hFFFFFFE2,
		32'h0000022B,
		32'h0000008D,
		32'h0000008C,
		32'hFFFFFED4,
		32'hFFFFFBF7,
		32'hFFFFFF23,
		32'h00000494,
		32'h00000110,
		32'h00000103,
		32'hFFFFFE51,
		32'h000003C7,
		32'h000003BD,
		32'h00000134,
		32'h000003FA,
		32'h0000006F,
		32'h0000001D,
		32'h0000018B,
		32'hFFFFFA98,
		32'h00000396,
		32'hFFFFFD12,
		32'hFFFFFD8D,
		32'hFFFFFFAB,
		32'hFFFFFBC6,
		32'hFFFFFC62,
		32'h0000048C,
		32'hFFFFFF15,
		32'h0000020F,
		32'h0000011F,
		32'h00000583,
		32'hFFFFFD5D,
		32'hFFFFFD1F,
		32'h00000562,
		32'hFFFFFC41,
		32'hFFFFFA78,
		32'hFFFFFF03,
		32'h0000032E,
		32'h00000282,
		32'hFFFFFC3A,
		32'hFFFFFBA5,
		32'h000001CF,
		32'hFFFFFC51
	};
	assign bias[31:0] = mem[a1];
        assign bias[63:32] = mem[a2];
        assign bias[95:64] = mem[a3];
        assign bias[127:96] = mem[a4];
endmodule

