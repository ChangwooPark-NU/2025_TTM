`timescale 1ns/1ps 

module regfile1 ( 
	input logic clk, 
	input logic [6:0] a1, a2, a3, a4,
	output logic [127:0] bias
); 
	logic [31:0] mem [0:127] = '{ 
		32'h00000082,
		32'hFFFFFA8C,
		32'hFFFFFE90,
		32'hFFFFFF81,
		32'h00000419,
		32'h000003B0,
		32'hFFFFFCE6,
		32'h000002A2,
		32'h00000114,
		32'hFFFFFC7A,
		32'hFFFFFDDE,
		32'h00000139,
		32'h0000027C,
		32'hFFFFFE23,
		32'h000001B8,
		32'h000000D6,
		32'hFFFFFB55,
		32'hFFFFFF79,
		32'h00000173,
		32'h000001D2,
		32'h0000003A,
		32'hFFFFFCFE,
		32'hFFFFFE67,
		32'h000002F2,
		32'h0000034D,
		32'hFFFFFFED,
		32'h0000064B,
		32'h0000017D,
		32'hFFFFFBFC,
		32'h00000005,
		32'hFFFFFF6E,
		32'h0000000B,
		32'h0000019A,
		32'hFFFFFF5E,
		32'hFFFFFCE8,
		32'h000003AD,
		32'h00000317,
		32'hFFFFFCCE,
		32'hFFFFFF1D,
		32'h00000294,
		32'hFFFFFF5C,
		32'h000000EA,
		32'hFFFFFD89,
		32'hFFFFFD90,
		32'hFFFFFB8B,
		32'h0000063D,
		32'h000004FA,
		32'h0000048C,
		32'hFFFFFF0D,
		32'hFFFFFE05,
		32'h00000245,
		32'h00000351,
		32'hFFFFFFEA,
		32'hFFFFFF1E,
		32'hFFFFF9BA,
		32'hFFFFFCA3,
		32'h0000010F,
		32'h0000000D,
		32'h000000CF,
		32'h000004FA,
		32'h00000359,
		32'hFFFFFBC4,
		32'hFFFFFAA3,
		32'h000000B4,
		32'h000002DA,
		32'hFFFFFADA,
		32'h0000022C,
		32'hFFFFFC80,
		32'h000002CB,
		32'hFFFFFD8A,
		32'h00000552,
		32'h000004A8,
		32'hFFFFFCAD,
		32'hFFFFFB26,
		32'h000001E2,
		32'h00000449,
		32'h0000029F,
		32'hFFFFFD3A,
		32'h000004DD,
		32'hFFFFFB12,
		32'h000004B5,
		32'hFFFFFD8F,
		32'hFFFFFF91,
		32'hFFFFFF9D,
		32'hFFFFFDF0,
		32'hFFFFFEC6,
		32'h00000200,
		32'h00000101,
		32'h000000CE,
		32'h00000621,
		32'hFFFFFFEF,
		32'hFFFFFC80,
		32'hFFFFFA11,
		32'h00000555,
		32'hFFFFFBCF,
		32'h00000141,
		32'hFFFFFCC5,
		32'hFFFFFC55,
		32'h00000163,
		32'h00000441,
		32'hFFFFF9FC,
		32'h0000001B,
		32'hFFFFFCB5,
		32'h000000B5,
		32'hFFFFFD74,
		32'hFFFFF9B0,
		32'hFFFFFB41,
		32'hFFFFFD5C,
		32'hFFFFFBA9,
		32'h00000099,
		32'hFFFFFD7F,
		32'hFFFFFD89,
		32'hFFFFFDEC,
		32'h0000024C,
		32'hFFFFFEB5,
		32'h0000057F,
		32'h000001F3,
		32'hFFFFFA15,
		32'hFFFFFFA4,
		32'hFFFFFA35,
		32'h00000334,
		32'hFFFFFD1A,
		32'h0000007E,
		32'h00000238,
		32'h00000790,
		32'hFFFFFF4E,
		32'hFFFFFFE9,
		32'h000004CA
        }; 	
	assign bias[31:0] = mem[a1]; 
	assign bias[63:32] = mem[a2]; 
	assign bias[95:64] = mem[a3]; 
	assign bias[127:96] = mem[a4]; 
endmodule 


