`timescale 1ns/1ps 

module regfile3 ( 
	input logic clk, 
	input logic [6:0] a1, a2, a3, a4,
	output logic [127:0] bias
); 
	logic [31:0] mem [0:127] = '{ 
		32'hFFFFF9F5,
		32'hFFFFFB35,
		32'hFFFFFD60,
		32'h0000033C,
		32'h000003A0,
		32'h00000306,
		32'h0000027B,
		32'h00000440,
		32'h00000289,
		32'hFFFFFD31,
		32'hFFFFFCB7,
		32'h000003F7,
		32'hFFFFFE37,
		32'hFFFFFD12,
		32'h000000EC,
		32'hFFFFFBEC,
		32'h00000046,
		32'h000006EC,
		32'h00000382,
		32'hFFFFFEE4,
		32'h00000149,
		32'h00000241,
		32'hFFFFFCD9,
		32'hFFFFFE5F,
		32'h00000483,
		32'hFFFFFC31,
		32'h000002AD,
		32'hFFFFFC78,
		32'h00000102,
		32'hFFFFFDA1,
		32'h00000421,
		32'hFFFFFCD5,
		32'hFFFFFCA3,
		32'h00000337,
		32'hFFFFFF40,
		32'h00000623,
		32'hFFFFFC65,
		32'h0000050F,
		32'h0000010A,
		32'h0000057A,
		32'hFFFFFF4A,
		32'hFFFFFDA2,
		32'h0000002D,
		32'hFFFFFC60,
		32'hFFFFFFE4,
		32'hFFFFFB3F,
		32'h0000040A,
		32'h000005E7,
		32'hFFFFFED0,
		32'h00000061,
		32'h00000296,
		32'hFFFFFF7E,
		32'hFFFFFEAD,
		32'hFFFFFD45,
		32'h000005D9,
		32'h00000074,
		32'h000004D7,
		32'h00000522,
		32'h00000537,
		32'hFFFFFF5C,
		32'hFFFFFE88,
		32'hFFFFFDD4,
		32'h00000748,
		32'hFFFFFCDA,
		32'hFFFFFFA2,
		32'hFFFFFBB5,
		32'hFFFFF85F,
		32'hFFFFFFD6,
		32'hFFFFFCFE,
		32'hFFFFFA9E,
		32'hFFFFFE94,
		32'h000005F4,
		32'h000000A5,
		32'h00000173,
		32'hFFFFFB62,
		32'hFFFFFDA2,
		32'h00000472,
		32'h000005A2,
		32'hFFFFFED8,
		32'hFFFFFC5C,
		32'h000006FB,
		32'hFFFFFCDE,
		32'hFFFFFC27,
		32'h000002F3,
		32'hFFFFFFF5,
		32'hFFFFFFFA,
		32'h0000035E,
		32'h00000420,
		32'h0000066E,
		32'h00000475,
		32'h00000051,
		32'h000004BD,
		32'hFFFFF8D3,
		32'hFFFFFD9E,
		32'hFFFFFA03,
		32'hFFFFFD89,
		32'h000003FF,
		32'hFFFFFFEF,
		32'hFFFFFD95,
		32'h00000027,
		32'hFFFFFD5B,
		32'hFFFFFFE0,
		32'h00000556,
		32'hFFFFFB06,
		32'h000002AD,
		32'h00000169,
		32'h000005A6,
		32'hFFFFFE18,
		32'hFFFFFEE9,
		32'hFFFFFD8C,
		32'hFFFFFF94,
		32'hFFFFFAB2,
		32'hFFFFFBFF,
		32'h0000016C,
		32'hFFFFFF8E,
		32'h0000039C,
		32'h0000006B,
		32'hFFFFFCDC,
		32'hFFFFFA04,
		32'hFFFFFAC4,
		32'h0000009C,
		32'hFFFFFF99,
		32'h00000543,
		32'h00000678,
		32'h000005D5,
		32'h00000379,
		32'h00000569,
		32'hFFFFFECE
	}; 
	assign bias[31:0] = mem[a1];
        assign bias[63:32] = mem[a2];
        assign bias[95:64] = mem[a3];
        assign bias[127:96] = mem[a4];
endmodule

